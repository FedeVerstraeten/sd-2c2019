package parametersPackage is
    constant NCOBITS : integer :=  12;
    constant FREQCONTROLBITS : integer := 11;
    constant DATABITS : integer := 8;
end parametersPackage;
